package version is
    constant GIT_VERSION : natural := 16#73400cd#;
    constant GIT_DIRTY : natural := 1;
    constant VERSION_MAJOR : natural := 0;
    constant VERSION_MINOR : natural := 1;
    constant VERSION_PATCH : natural := 0;
end;
