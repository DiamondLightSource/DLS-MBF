-- Sequential state machine to compute angle and magnitude of vector iq_i.
-- Processing is initiated by pulsing start_i and completion signalled by
-- done_o.
--
-- The algorithm implemented here is the classic CORDIC algorithm:
--
--      Volder, J.E., 1959; "The CORDIC Trigonometric Computing Technique",
--      IRE Transactions on Electronic Computers, V.  EC-8, No. 3, pp. 330-334
--
-- The basic iteration step is the calculation:
--
--      x <= x + (y >>> n)
--      y <= y - (x >>> n)
--
-- which can be written as (let xy = column vector of x and y):
--
--            [1    2^-n]
--      xy <= [-2^-n   1] xy = sqrt(1 + 2^-2n) R(th) xy , where tan(th) = 2^-n
--
-- where R(th) is the rotation matrix to rotate a vectory by angle th, in this
-- case tan^-1(2^-n).  Here we perform a sequence of positive or negative
-- rotations for increasing values of n to drive one component of the vector to
-- zero.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.defines.all;
use work.support.all;

use work.nco_defs.all;

entity tune_pll_cordic is
    port (
        clk_i : in std_ulogic;

        iq_i : in cos_sin_t;
        start_i : in std_ulogic;

        angle_o : out signed;
        magnitude_o : out unsigned;
        done_o : out std_ulogic := '0'
    );
end;

architecture arch of tune_pll_cordic is
    -- The number of available angle bits is determined by the autogenerated
    -- cordic_table entity
    constant ANGLE_BITS : natural := 18;
    -- The top two bits of the computed angle are derived directly from the
    -- quadrant, the rest will need to be shifted in
    constant SHIFT_COUNT : natural := ANGLE_BITS - 2;
    -- This word size includes two extra low-order bits for rounding included in
    -- the arc-tangent result
    constant ROUNDING_BITS : natural := 2;
    constant ATAN_BITS : natural := ANGLE_BITS + ROUNDING_BITS;

    constant WORD_SIZE_IN : natural := iq_i.cos'LENGTH;
    constant MAX_NORMALISE_SHIFT : natural := 15;

    -- To account for CORDIC growth, a factor of around 1.65 together with a
    -- further factor of sqrt(2) from rotation, we need two more bits of high
    -- order result.  We'll return this entire result as the magnitude.
    constant IQ_SIZE : natural := magnitude_o'LENGTH + 2;


    -- Inverse tangent
    subtype cordic_angle_t is signed(ATAN_BITS-1 downto 0);
    signal atan : cordic_angle_t;
    signal angle_update : cordic_angle_t;

    -- Cordic state machine.
    type state_t is (STATE_IDLE, STATE_NORMALISE, STATE_SHIFT, STATE_ADD);
    signal state : state_t := STATE_IDLE;
    signal step_count : unsigned(bits(SHIFT_COUNT-1)-1 downto 0)
        := (others => '0');
    signal done : std_ulogic := '0';

    signal quadrant : std_ulogic_vector(1 downto 0);

    signal normalised : boolean;
    signal normalise_shift : unsigned(bits(MAX_NORMALISE_SHIFT)-1 downto 0);
    signal iq_normal : iq_i'SUBTYPE;

    subtype iq_accum_t is cos_sin_t(
        cos(IQ_SIZE-1 downto 0), sin(IQ_SIZE-1 downto 0));

    signal iq : iq_accum_t;
    signal shifted : iq_accum_t;
    signal angle : signed(ATAN_BITS-1 downto 0);


    function initial_angle(quadrant : integer) return cordic_angle_t is
    begin
        return to_signed(quadrant, 2) & to_signed(0, ATAN_BITS - 2);
    end;

begin
    assert angle_o'LENGTH = ANGLE_BITS severity failure;

    -- Angle adustment for step lookup.
    atan_table : entity work.cordic_table port map (
        addr_i => step_count,
        dat_o => atan
    );

    quadrant <= sign_bit(iq_i.cos) & sign_bit(iq_i.sin);

    normalised <=
        normalise_shift = MAX_NORMALISE_SHIFT or
        iq_normal.cos(WORD_SIZE_IN-2) = '1' or
        iq_normal.sin(WORD_SIZE_IN-2) = '1';

    process (clk_i) begin
        if rising_edge(clk_i) then
            -- Cordic state machine
            case state is
                when STATE_IDLE =>
                    done <= '0';
                    step_count <= (others => '0');
                    normalise_shift <= (others => '0');
                    if start_i = '1' then
                        state <= STATE_NORMALISE;
                    end if;

                    -- For the first rotation rotate into first quadrant so both
                    -- components are non-negative
                    case quadrant is
                        -- Note that we use complement rather than negation to
                        -- avoid a rather gratuitous extra bit of growth (for
                        -- min_int), at the cost of 1 bottom bit error.
                        when "00" =>    -- 0 deg rotation
                            iq_normal.cos <= iq_i.cos;
                            iq_normal.sin <= iq_i.sin;
                            angle <= initial_angle(0);
                        when "10" =>    -- 90 deg rotation
                            iq_normal.cos <= iq_i.sin;
                            iq_normal.sin <= not iq_i.cos;
                            angle <= initial_angle(1);
                        when "11" =>    -- 180 deg rotation
                            iq_normal.cos <= not iq_i.cos;
                            iq_normal.sin <= not iq_i.sin;
                            angle <= initial_angle(-2);
                        when "01" =>    -- 270 deg rotation
                            iq_normal.cos <= not iq_i.sin;
                            iq_normal.sin <= iq_i.cos;
                            angle <= initial_angle(-1);
                        when others =>
                    end case;

                when STATE_NORMALISE =>
                    if normalised then
                        -- Value is already normalised, move on to next step
                        iq.cos <= "00" & iq_normal.cos;
                        iq.sin <= "00" & iq_normal.sin;
                        state <= STATE_SHIFT;
                    else
                        -- Shift and go around
                        iq_normal.cos <= shift_left(iq_normal.cos, 1);
                        iq_normal.sin <= shift_left(iq_normal.sin, 1);
                        normalise_shift <= normalise_shift + 1;
                    end if;


                when STATE_SHIFT =>
                    state <= STATE_ADD;
                    shifted.cos <= shift_right(iq.cos, to_integer(step_count));
                    shifted.sin <= shift_right(iq.sin, to_integer(step_count));
                    angle_update <= atan;

                when STATE_ADD =>
                    if step_count = SHIFT_COUNT - 1 then
                        done <= '1';
                        state <= STATE_IDLE;
                    else
                        step_count <= step_count + 1;
                        state <= STATE_SHIFT;
                    end if;

                    if iq.sin >= 0 then
                        iq.cos <= iq.cos + shifted.sin;
                        iq.sin <= iq.sin - shifted.cos;
                        angle <= angle + angle_update;
                    else
                        iq.cos <= iq.cos - shifted.sin;
                        iq.sin <= iq.sin + shifted.cos;
                        angle <= angle - angle_update;
                    end if;
            end case;

            -- Register the final result
            if done = '1' then
                -- Discard the sign bit for our unsigned result
                magnitude_o <= shift_right(unsigned(
                    iq.cos(IQ_SIZE-2 downto IQ_SIZE - magnitude_o'LENGTH-1)),
                    to_integer(normalise_shift));
                angle_o <= angle(ATAN_BITS-1 downto ROUNDING_BITS);
            end if;
            done_o <= done;
        end if;
    end process;
end;
