library ieee;
use ieee.std_logic_1164.all;

entity interconnect_wrapper is
    port (
        C0_DDR3_addr : out std_logic_vector(14 downto 0);
        C0_DDR3_ba : out std_logic_vector(2 downto 0);
        C0_DDR3_cas_n : out std_logic;
        C0_DDR3_ck_n : out std_logic_vector(0 to 0);
        C0_DDR3_ck_p : out std_logic_vector(0 to 0);
        C0_DDR3_cke : out std_logic_vector(0 to 0);
        C0_DDR3_dm : out std_logic_vector(7 downto 0);
        C0_DDR3_dq : inout std_logic_vector(63 downto 0);
        C0_DDR3_dqs_n : inout std_logic_vector(7 downto 0);
        C0_DDR3_dqs_p : inout std_logic_vector(7 downto 0);
        C0_DDR3_odt : out std_logic_vector(0 to 0);
        C0_DDR3_ras_n : out std_logic;
        C0_DDR3_reset_n : out std_logic;
        C0_DDR3_we_n : out std_logic;
        C1_DDR3_addr : out std_logic_vector(12 downto 0);
        C1_DDR3_ba : out std_logic_vector(2 downto 0);
        C1_DDR3_cas_n : out std_logic;
        C1_DDR3_ck_n : out std_logic_vector(0 to 0);
        C1_DDR3_ck_p : out std_logic_vector(0 to 0);
        C1_DDR3_cke : out std_logic_vector(0 to 0);
        C1_DDR3_dm : out std_logic_vector(1 downto 0);
        C1_DDR3_dq : inout std_logic_vector(15 downto 0);
        C1_DDR3_dqs_n : inout std_logic_vector(1 downto 0);
        C1_DDR3_dqs_p : inout std_logic_vector(1 downto 0);
        C1_DDR3_odt : out std_logic_vector(0 to 0);
        C1_DDR3_ras_n : out std_logic;
        C1_DDR3_reset_n : out std_logic;
        C1_DDR3_we_n : out std_logic;
        CLK200MHZ : in std_logic;
        CLK533MHZ0_clk_n : in std_logic;
        CLK533MHZ0_clk_p : in std_logic;
        CLK533MHZ1_clk_n : in std_logic;
        CLK533MHZ1_clk_p : in std_logic;
        DSP_CLK : in std_logic;
        DSP_RESETN : in std_logic;
        FCLKA : in std_logic;
        INTR : in std_logic_vector(30 downto 0);
        M_DSP_REGS_araddr : out std_logic_vector(15 downto 0);
        M_DSP_REGS_arprot : out std_logic_vector(2 downto 0);
        M_DSP_REGS_arready : in std_logic;
        M_DSP_REGS_arvalid : out std_logic;
        M_DSP_REGS_awaddr : out std_logic_vector(15 downto 0);
        M_DSP_REGS_awprot : out std_logic_vector(2 downto 0);
        M_DSP_REGS_awready : in std_logic;
        M_DSP_REGS_awvalid : out std_logic;
        M_DSP_REGS_bready : out std_logic;
        M_DSP_REGS_bresp : in std_logic_vector(1 downto 0);
        M_DSP_REGS_bvalid : in std_logic;
        M_DSP_REGS_rdata : in std_logic_vector(31 downto 0);
        M_DSP_REGS_rready : out std_logic;
        M_DSP_REGS_rresp : in std_logic_vector(1 downto 0);
        M_DSP_REGS_rvalid : in std_logic;
        M_DSP_REGS_wdata : out std_logic_vector(31 downto 0);
        M_DSP_REGS_wready : in std_logic;
        M_DSP_REGS_wstrb : out std_logic_vector(3 downto 0);
        M_DSP_REGS_wvalid : out std_logic;
        REG_CLK : in std_logic;
        REG_RESETN : in std_logic;
        S_DSP_DRAM0_awaddr : in std_logic_vector(47 downto 0);
        S_DSP_DRAM0_awburst : in std_logic_vector(1 downto 0);
        S_DSP_DRAM0_awcache : in std_logic_vector(3 downto 0);
        S_DSP_DRAM0_awlen : in std_logic_vector(7 downto 0);
        S_DSP_DRAM0_awlock : in std_logic_vector(0 to 0);
        S_DSP_DRAM0_awprot : in std_logic_vector(2 downto 0);
        S_DSP_DRAM0_awqos : in std_logic_vector(3 downto 0);
        S_DSP_DRAM0_awready : out std_logic;
        S_DSP_DRAM0_awregion : in std_logic_vector(3 downto 0);
        S_DSP_DRAM0_awsize : in std_logic_vector(2 downto 0);
        S_DSP_DRAM0_awvalid : in std_logic;
        S_DSP_DRAM0_bready : in std_logic;
        S_DSP_DRAM0_bresp : out std_logic_vector(1 downto 0);
        S_DSP_DRAM0_bvalid : out std_logic;
        S_DSP_DRAM0_wdata : in std_logic_vector(63 downto 0);
        S_DSP_DRAM0_wlast : in std_logic;
        S_DSP_DRAM0_wready : out std_logic;
        S_DSP_DRAM0_wstrb : in std_logic_vector(7 downto 0);
        S_DSP_DRAM0_wvalid : in std_logic;
        S_DSP_DRAM1_awaddr : in std_logic_vector(47 downto 0);
        S_DSP_DRAM1_awprot : in std_logic_vector(2 downto 0);
        S_DSP_DRAM1_awready : out std_logic;
        S_DSP_DRAM1_awvalid : in std_logic;
        S_DSP_DRAM1_bready : in std_logic;
        S_DSP_DRAM1_bresp : out std_logic_vector(1 downto 0);
        S_DSP_DRAM1_bvalid : out std_logic;
        S_DSP_DRAM1_wdata : in std_logic_vector(63 downto 0);
        S_DSP_DRAM1_wready : out std_logic;
        S_DSP_DRAM1_wstrb : in std_logic_vector(7 downto 0);
        S_DSP_DRAM1_wvalid : in std_logic;
        nCOLDRST : in std_logic;
        pcie_mgt_rxn : in std_logic_vector(7 downto 0);
        pcie_mgt_rxp : in std_logic_vector(7 downto 0);
        pcie_mgt_txn : out std_logic_vector(7 downto 0);
        pcie_mgt_txp : out std_logic_vector(7 downto 0)
   );
end;

architecture arch of interconnect_wrapper is
begin
end;
